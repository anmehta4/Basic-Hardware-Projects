module ALU_tb();

  //////////////////////////////////
  // Define stimulus of type reg //
  ////////////////////////////////
  reg [7:0] A,B;
  reg [1:0] mode;
  reg error;	// set if an error occurred during testing
  
  ////////////////////////////////////////////////////
  // Signals hooked to DUT output are of type wire //
  //////////////////////////////////////////////////
  wire [7:0] result;
  
  //////////////////////
  // Instantiate DUT //
  ////////////////////
  ALU iDUT(.A(A), .B(B), .mode(mode), .Y(result));
  
  initial begin
    error = 0;		// innocent till proven guilty
	
	$display("Performing mode 00 testing");
    mode = 2'b00;	// start testing Shift Right Arithmetic
	A = 8'hAA;
	B = 8'h56;
	#1;
	if (result!==8'h2B) begin
	  $display("ERR: SRA(0x56) should result in 0x2B.  Your answer was %h",result);
	  error = 1;
	end
	
	B = 8'hAB;
	#1;
	if (result!==8'hD5) begin
	  $display("ERR: SRA(0xAB) should result in 0xD5.  Your answer was %h",result);
	  error = 1;
	end
	
	if (!error)
	  $display("Good...you passed mode 00 moving to mode 01 next");
	  
	mode = 2'b01;
	B = 8'h6E;
	#1;
	if (result!==8'hDC) begin
	  $display("ERR: 0x6E*2 should result in 0xDC.  Your answer was %h",result);
	  error = 1;
	end	else
	  $display("Good...you passed mode 01 moving to mode 10 next");
	  
	mode = 2'b10;
	A = 8'h95;
	#1;
	if (result!==8'h03) begin
	  $display("ERR: 0x95 + 0x6E should result in 0x03.  Your answer was %h",result);
	  error = 1;
	end	
	B = 8'h4A;
	#1;
	if (result!==8'hDF) begin
	  $display("ERR: 0x95 + 0x4A should result in 0xDF.  Your answer was %h",result);
	  error = 1;
	end

	if (!error)
	  $display("Good...you passed mode 10 moving to mode 11 next");
	  
	mode = 2'b11;
	A = 8'h9C;
	#1;
	if (result!==8'h52) begin
	  $display("ERR: 0x9C - 0x4A should result in 0x52.  Your answer was %h",result);
	  error = 1;
	end	
	A = 8'h56;
	B = 8'h7D;
	#1;
	if (result!==8'hD9) begin
	  $display("ERR: 0x56 - 0x7D should result in 0xD9.  Your answer was %h",result);
	  error = 1;
	end	

    if (!error)
      $display("YAHOO!! test passed");
    
    $stop();
	
  end
  
endmodule
